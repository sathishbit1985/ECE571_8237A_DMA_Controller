////////////////////////////////////////////////////////////////////////////////////
//////--------- ECE571_SPRING2022 FINAL PROJECT ------------------------------
/////---------- DMA CONTROLLER ---------------------------------------------
/////---------- TEST BENCH FOR VERIFICATION -------------------------------  
/////----------- VERIFICATION TEAM MEMBERS: Manoj, Kaavya, Saket -------------
//////////////////////////////////////////////////////////////////////////////////

module top();
  
  
endmodule
